module adder(input [31:0] A, B, output [31:0] adder_out);
	
	assign adder_out = A + B;	

endmodule
